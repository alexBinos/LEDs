

module pwm_generator #(
   parameter integer SYS_CLK_FREQ = 100_000_000
)(
   input wire clk_in,
   input wire n_reset_in,
   input wire [7:0]
);

endmodule
