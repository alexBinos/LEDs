

module led_display_pattern_gen #(
   parameter integer SYS_CLK_FREQ = 100_000_000
)(
   input  wire clk_in,
   input  wire n_reset_in
);
   
endmodule
